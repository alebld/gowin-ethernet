module mdio (
	     input porco
	     );
   input ret;
   
   
   
